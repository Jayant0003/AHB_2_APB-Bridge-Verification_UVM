class apb_slave_agent extends uvm_agent;
`uvm_component_utils(apb_slave_agent)


apb_slave_agent_config apb_agent_cfg;
apb_slave_driver drvh;
apb_slave_monitor monh;
apb_slave_sequencer seqrh;
function new(string name=get_type_name(),uvm_component parent);
	super.new(name,parent);
endfunction

function void build_phase(uvm_phase phase);
	super.build_phase(phase);
	if(!uvm_config_db #(apb_slave_agent_config)::get(this,"","apb_slave_agent_config",apb_agent_cfg))
	`uvm_fatal(get_type_name,"error while getting agent_cfg");

	monh=apb_slave_monitor::type_id::create("monh",this);
	if(apb_agent_cfg.is_active==UVM_ACTIVE) begin
	drvh=apb_slave_driver::type_id::create("drvh",this);
	seqrh=apb_slave_sequencer::type_id::create("seqrh",this);
	end
	
		
endfunction
function void connect_phase(uvm_phase phase);
	super.connect_phase(phase);
	drvh.seq_item_port.connect(seqrh.seq_item_export);
endfunction

endclass

