package test_pkg;
import uvm_pkg::*;
`include "definitions.v"
`include "uvm_macros.svh"
`include "ahb_master_agent_config.sv"
`include "apb_slave_agent_config.sv"
`include "env_config.sv"

`include "slave_xtn.sv"
`include "slave_seqs.sv"
`include "apb_slave_sequencer.sv"
`include "apb_slave_driver.sv"
`include "apb_slave_monitor.sv"
`include "apb_slave_agent.sv"
`include "apb_slave_agent_top.sv"


`include "master_xtn.sv"
`include "master_seqs.sv"
`include "ahb_master_sequencer.sv"
`include "ahb_master_driver.sv"
`include "ahb_master_monitor.sv"
`include "ahb_master_agent.sv"
`include "ahb_master_agent_top.sv"


`include "scoreboard.sv"
`include "virtual_sequencer.sv"
`include "virtual_seqs.sv"
`include "tb.sv"

`include "test_lib.sv"
endpackage
