class slave_seqs extends uvm_sequence#(slave_xtn);
`uvm_object_utils(slave_seqs)

function new(string name=get_type_name);
	super.new(name);
endfunction


endclass
